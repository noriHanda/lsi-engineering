module rom_10bit_64word(AD,
                        Q);
    input [5:0] AD;
    output [9:0] Q;
    
    reg [9:0] q [0:63];
    
    initial begin
        // Hazardous code
        // q[6'd0]  <= {4'b0111, 6'd63};
        // q[6'd1]  <= {4'b1100, 6'd0};
        // q[6'd2]  <= {4'b0110, 6'd1};
        // q[6'd3]  <= {4'b0001, 6'd1};
        // q[6'd4]  <= {4'b0110, 6'd1};
        // q[6'd5]  <= {4'b1100, 6'd3};
        // q[6'd6]  <= {4'b0111, 6'd63};
        // q[6'd7]  <= {4'b1100, 6'd6};
        // q[6'd8]  <= {4'b0110, 6'd1};
        // q[6'd9]  <= {4'b0110, 6'd1};
        // q[6'd10] <= {4'b0001, 6'd1};
        // q[6'd11] <= {4'b1100, 6'd9};
        // q[6'd12] <= {4'b1001, 6'd0};
        // q[6'd13] <= {4'b1011, 6'd13};
        
        // Fixed code
        q[6'd0]  <= {4'b0111, 6'd63};
        q[6'd1]  <= {4'b1100, 6'd0 };
        q[6'd2]  <= {4'b0000, 6'd0 };
        q[6'd3]  <= {4'b0000, 6'd0 };
        q[6'd4]  <= {4'b0000, 6'd0 };
        q[6'd5]  <= {4'b0110, 6'd1 };
        q[6'd6]  <= {4'b0001, 6'd1 };
        q[6'd7]  <= {4'b0110, 6'd1 };
        q[6'd8]  <= {4'b1100, 6'd6 };
        q[6'd9]  <= {4'b0000, 6'd0 };
        q[6'd10] <= {4'b0000, 6'd0 };
        q[6'd11] <= {4'b0000, 6'd0 };
        q[6'd12] <= {4'b0111, 6'd63};
        q[6'd13] <= {4'b1100, 6'd12};
        q[6'd14] <= {4'b0000, 6'd0 };
        q[6'd15] <= {4'b0000, 6'd0 };
        q[6'd16] <= {4'b0000, 6'd0 };
        q[6'd17] <= {4'b0110, 6'd1 };
        q[6'd18] <= {4'b0000, 6'd0 };
        q[6'd19] <= {4'b0110, 6'd1 };
        q[6'd20] <= {4'b0001, 6'd1 };
        q[6'd21] <= {4'b1100, 6'd19};
        q[6'd22] <= {4'b0000, 6'd0 };
        q[6'd23] <= {4'b0000, 6'd0 };
        q[6'd24] <= {4'b0000, 6'd0 };
        q[6'd25] <= {4'b1001, 6'd0 };
        q[6'd26] <= {4'b1011, 6'd26};
        q[6'd27] <= {4'b0000, 6'd0 };
        q[6'd28] <= {4'b0000, 6'd0 };
        q[6'd29] <= {4'b0000, 6'd0 };
    end
    
    assign Q = q[AD];
endmodule
