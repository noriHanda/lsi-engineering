`include "dec_7seg.v"

module accumulator(CLK, RST_N, B, LEDB, LEDC, HEXB1, HEXB0, HEXA1, HEXA0);
	input CLK;// 50MHz
	input RST_N;
	input [3:0] B;
	output [3:0] LEDB;
	output LEDC;
	output [6:0] HEXB1, HEXB0, HEXA1, HEXA0;

	// Please write down your code!



endmodule