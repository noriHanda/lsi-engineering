`include "dec_7seg.v"

module shift_reg(CLK, RST_N, D, LEDD, LEDC, HEXq7, HEXq6, HEXq5, HEXq4, HEXq3, HEXq2, HEXq1, HEXq0);
	input CLK;// 50MHz
	input RST_N;
	input [3:0] D;
	output [3:0] LEDD;
	output LEDC;
	output [6:0] HEXq7, HEXq6, HEXq5, HEXq4, HEXq3, HEXq2, HEXq1, HEXq0;

	// Please write down your code!



endmodule