module rom_10bit_64word(AD,
                        Q);
    input [5:0] AD;
    output [9:0] Q;
    
    reg [9:0] q [0:63];
    
    initial begin
        // 課題1 (#12 P18) のプログラム
        // q[6'd0] <= {4'b0100, 6'd5};// MOV A, 5
        // q[6'd1] <= {4'b1000, 6'd10};// MOV B, 10
        
        // 課題2 (#12 P21) のプログラム
        // q[6'd0] <= {4'b0100, 6'd5};// MOV A, 5
        // q[6'd1] <= {4'b0000, 6'd0};// NOP
        // q[6'd2] <= {4'b0001, 6'd1};// NOP
        
        // 課題3 (#12 P25) のプログラム
        // q[6'd0] <= {4'b1011, 6'd5};
        // q[6'd1] <= {4'b0000, 6'd0};
        // q[6'd2] <= {4'b0000, 6'd0};
        // q[6'd3] <= {4'b0000, 6'd0};
        // q[6'd4] <= {4'b0100, 6'd4};
        // q[6'd5] <= {4'b1010, 6'd1};
        
        // 課題4 (#12 P26) のプログラム
        q[6'd0] <= {4'b0100, 6'd62};
        q[6'd1] <= {4'b0000, 6'd0};
        q[6'd2] <= {4'b0001, 6'd1};
        q[6'd3] <= {4'b1100, 6'd2};
        q[6'd4] <= {4'b0000, 6'd0};
        q[6'd5] <= {4'b0000, 6'd0};
        q[6'd6] <= {4'b0000, 6'd0};
    end
    
    assign Q = q[AD];
endmodule
