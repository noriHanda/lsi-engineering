module x_scan (
    input x0, x1, x2,
);

endmodule // x_scan

module y_scan (
    
);

endmodule // y_scan