`include "dec_7seg.v"

module adder(A, B, LEDA, LEDB, LEDY, HEXA, HEXB, HEXY);
	input [2:0] A, B;
	output [2:0] LEDA, LEDB;
	output [3:0] LEDY;
	output [6:0] HEXA, HEXB, HEXY;

	wire [3:0] Y;

	// Please write down your code!



endmodule