module led_flash(CLK, RST_N, LED);
	input CLK;// 50MHz
	input RST_N;
	output LED;

	reg LED_025Hz;// 0.25Hz

	// Please write down your code!



endmodule