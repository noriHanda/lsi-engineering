module DataSource (
    
);

endmodule //DataSource