`include "dec_7seg.v"

module comparator(A, B, LEDA, LEDB, HEXA, HEXB, HEXC);
	input [3:0] A, B;
	output [3:0] LEDA, LEDB;
	output [6:0] HEXA, HEXB, HEXC;

	// Please write down your code!



endmodule